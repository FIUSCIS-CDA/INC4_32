///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: INC4_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: A (32-bit)
reg[31:0] A;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Outputs: S (32-bit)
wire[31:0] S;
///////////////////////////////////////////////////////////////////////////////////

INC4_32 myAdder(.A(A), .S(S));

initial begin
/////////////////////////////////////////////////////////////////////////////
// Test: A=45
$display("Testing A=45: ");
A=45;  #10; 
verifyEqual32(S, A+4);
/////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end


endmodule